// This Verilog file automatically generated from controller.asm
//
module serial_wb_program(clk_i, pm_addr_i, pm_insn_o);
   input         clk_i;
   input  [9:0]  pm_addr_i;
   output [15:0] pm_insn_o;

   wire          clk_i;
   wire [9:0]    pm_addr_i;
   reg  [15:0]   pm_insn_o;



   always @(posedge clk_i)
       case(pm_addr_i)
        10'h000: pm_insn_o <= 16'h4f00; // 	set	#0x0,r15
        10'h001: pm_insn_o <= 16'hffff; // 	nop
        10'h002: pm_insn_o <= 16'hffff; // 	nop
        10'h003: pm_insn_o <= 16'h4000; // 	set	#0x0,r0
        10'h004: pm_insn_o <= 16'h4100; // 	set	#0x0,r1
        10'h005: pm_insn_o <= 16'h40ff; // 	set	#0xff,r0
        10'h006: pm_insn_o <= 16'h41ff; // 	set	#0xff,r1
        10'h007: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h008: pm_insn_o <= 16'h8407; // 	jmpc	delayloop
        10'h009: pm_insn_o <= 16'hffff; // 	nop
        10'h00a: pm_insn_o <= 16'h4040; // 	set	#0x40,r0
        10'h00b: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h00c: pm_insn_o <= 16'h4300; // 	set	LOW greetingstring,r3	; Pointer to greeting string
        10'h00d: pm_insn_o <= 16'h4405; // 	set	HIGH greetingstring,r4
        10'h00e: pm_insn_o <= 16'h87d3; // 	jsr	puts
        10'h00f: pm_insn_o <= 16'h400d; // 	set	#0x0d,r0	
        10'h010: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h011: pm_insn_o <= 16'h400a; // 	set	#0x0a,r0
        10'h012: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h013: pm_insn_o <= 16'h403e; // 	set	#0x3e,r0	; '>'
        10'h014: pm_insn_o <= 16'h8625; // 	jsr	putc		; print prompt
        10'h015: pm_insn_o <= 16'h8631; // 	jsr	getc		; get command character
        10'h016: pm_insn_o <= 16'h4144; // 	set	#0x44,r1	; 'D'
        10'h017: pm_insn_o <= 16'h1101; // 	xor	r0,r1,r1
        10'h018: pm_insn_o <= 16'h82cd; // 	jmpz	handle_logicanalyzer
        10'h019: pm_insn_o <= 16'hffff; // 	nop
        10'h01a: pm_insn_o <= 16'h4154; // 	set	#0x54,r1	;  'T' set trigger
        10'h01b: pm_insn_o <= 16'h1101; // 	xor	r0,r1,r1
        10'h01c: pm_insn_o <= 16'h8380; // 	jmpz	handle_settrigger
        10'h01d: pm_insn_o <= 16'hffff; // 	nop
        10'h01e: pm_insn_o <= 16'h4174; // 	set	#0x74,r1	;  't' trigger it
        10'h01f: pm_insn_o <= 16'h1101; // 	xor	r0,r1,r1
        10'h020: pm_insn_o <= 16'h8334; // 	jmpz	handle_trigger
        10'h021: pm_insn_o <= 16'hffff; // 	nop
        10'h022: pm_insn_o <= 16'h4007; // 	set	#0x7,r0		; ctrl g
        10'h023: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h024: pm_insn_o <= 16'h800f; // 	jmp	menuloop
        10'h025: pm_insn_o <= 16'h4101; // 	set	#0x1,r1
        10'h026: pm_insn_o <= 16'h9010; // 	out0	r1
        10'h027: pm_insn_o <= 16'h4202; // 	set	#0x2,r2		; UART_TX_IDLE
        10'h028: pm_insn_o <= 16'hffff; // 	nop
        10'h029: pm_insn_o <= 16'h5100; // 	in2	r1		; get status flags from UART
        10'h02a: pm_insn_o <= 16'h2112; // 	and	r1,r2,r1	; zero flag set if no TX slot available
        10'h02b: pm_insn_o <= 16'h8229; // 	jmpz	putc_waitidle
        10'h02c: pm_insn_o <= 16'hffff; // 	nop
        10'h02d: pm_insn_o <= 16'h4100; // 	set	#0x0,r1		; Output register of UART
        10'h02e: pm_insn_o <= 16'h9010; // 	out0	r1		; Address for TX transmit reg
        10'h02f: pm_insn_o <= 16'h9100; // 	out1	r0		; Transmit character
        10'h030: pm_insn_o <= 16'h8800; // 	rts
        10'h031: pm_insn_o <= 16'h4101; // 	set	#0x1,r1
        10'h032: pm_insn_o <= 16'h9010; // 	out0	r1
        10'h033: pm_insn_o <= 16'h4201; // 	set	#0x1,r2		; UART_RX_IDLE
        10'h034: pm_insn_o <= 16'hffff; // 	nop
        10'h035: pm_insn_o <= 16'h5100; // 	in2	r1
        10'h036: pm_insn_o <= 16'h2112; // 	and	r1,r2,r1
        10'h037: pm_insn_o <= 16'h8235; // 	jmpz	getc_waitchar
        10'h038: pm_insn_o <= 16'hffff; // 	nop
        10'h039: pm_insn_o <= 16'h4100; // 	set	#0x0,r1		; Address of RX recv reg
        10'h03a: pm_insn_o <= 16'h9010; // 	out0	r1
        10'h03b: pm_insn_o <= 16'hffff; // 	nop
        10'h03c: pm_insn_o <= 16'hffff; // 	nop
        10'h03d: pm_insn_o <= 16'h5000; // 	in2	r0		; Get character
        10'h03e: pm_insn_o <= 16'h4103; // 	set	#0x3,r1		; ctrl c
        10'h03f: pm_insn_o <= 16'h1101; // 	xor	r0,r1,r1
        10'h040: pm_insn_o <= 16'h8200; // 	jmpz	restart		; Restart if ctrl c was pressed
        10'h041: pm_insn_o <= 16'hffff; // 	nop
        10'h042: pm_insn_o <= 16'h8025; // 	jmp	putc		; Echo character
        10'h043: pm_insn_o <= 16'h4101; // 	set	#0x1,r1
        10'h044: pm_insn_o <= 16'h9010; // 	out0	r1
        10'h045: pm_insn_o <= 16'h4201; // 	set	#0x1,r2		; UART_RX_IDLE
        10'h046: pm_insn_o <= 16'hffff; // 	nop
        10'h047: pm_insn_o <= 16'h5100; // 	in2	r1
        10'h048: pm_insn_o <= 16'h2112; // 	and	r1,r2,r1
        10'h049: pm_insn_o <= 16'h8247; // 	jmpz	getc_quiet_waitchar
        10'h04a: pm_insn_o <= 16'hffff; // 	nop
        10'h04b: pm_insn_o <= 16'h4100; // 	set	#0x0,r1		; Address of RX recv reg
        10'h04c: pm_insn_o <= 16'h9010; // 	out0	r1
        10'h04d: pm_insn_o <= 16'hffff; // 	nop
        10'h04e: pm_insn_o <= 16'hffff; // 	nop
        10'h04f: pm_insn_o <= 16'h5000; // 	in2	r0		; Get character
        10'h050: pm_insn_o <= 16'h4103; // 	set	#0x3,r1		; ctrl c
        10'h051: pm_insn_o <= 16'h1101; // 	xor	r0,r1,r1
        10'h052: pm_insn_o <= 16'h8200; // 	jmpz	restart		; Restart if ctrl c was pressed
        10'h053: pm_insn_o <= 16'hffff; // 	nop
        10'h054: pm_insn_o <= 16'h8800; // 	rts
        10'h055: pm_insn_o <= 16'h4101; // 	set	#0x1,r1		; inc factor
        10'h056: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h057: pm_insn_o <= 16'h9140; // 	out1	r4
        10'h058: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h059: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h05a: pm_insn_o <= 16'h9150; // 	out1	r5
        10'h05b: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h05c: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h05d: pm_insn_o <= 16'h9160; // 	out1	r6
        10'h05e: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h05f: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h060: pm_insn_o <= 16'h9170; // 	out1	r7
        10'h061: pm_insn_o <= 16'h8800; // 	rts
        10'h062: pm_insn_o <= 16'h4101; // 	set	#0x01,r1	; increment constant
        10'h063: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h064: pm_insn_o <= 16'hffff; // 	nop			; Get rid of nop!
        10'h065: pm_insn_o <= 16'hffff; // 	nop
        10'h066: pm_insn_o <= 16'h5400; // 	in2	r4
        10'h067: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h068: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h069: pm_insn_o <= 16'hffff; // 	nop
        10'h06a: pm_insn_o <= 16'hffff; // 	nop
        10'h06b: pm_insn_o <= 16'h5500; // 	in2	r5
        10'h06c: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h06d: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h06e: pm_insn_o <= 16'hffff; // 	nop
        10'h06f: pm_insn_o <= 16'hffff; // 	nop
        10'h070: pm_insn_o <= 16'h5600; // 	in2	r6
        10'h071: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h072: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h073: pm_insn_o <= 16'hffff; // 	nop
        10'h074: pm_insn_o <= 16'hffff; // 	nop
        10'h075: pm_insn_o <= 16'h5700; // 	in2	r7
        10'h076: pm_insn_o <= 16'h8800; // 	rts
        10'h077: pm_insn_o <= 16'h8643; // 	jsr	getc_quiet
        10'h078: pm_insn_o <= 16'h41d0; // 	set	#0xd0,r1	; 0x100 - 0x30
        10'h079: pm_insn_o <= 16'h0101; // 	add	r0,r1,r1
        10'h07a: pm_insn_o <= 16'h847f; // 	jmpc	convascii_ge0	; jump if greater or equal to '0'
        10'h07b: pm_insn_o <= 16'hffff; // 	nop
        10'h07c: pm_insn_o <= 16'h4007; // 	set	#0x7,r0		; ctrl g
        10'h07d: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h07e: pm_insn_o <= 16'h8077; // 	jmp	getnibble	; restart nibbleloop
        10'h07f: pm_insn_o <= 16'h41c6; // 	set	#0xc6,r1	; 0x100 - 0x39
        10'h080: pm_insn_o <= 16'h0101; // 	add	r0,r1,r1
        10'h081: pm_insn_o <= 16'h8486; // 	jmpc	convascii_gt9
        10'h082: pm_insn_o <= 16'hffff; // 	nop
        10'h083: pm_insn_o <= 16'h41d0; // 	set	#0xd0,r1		; -0x30
        10'h084: pm_insn_o <= 16'h0301; // 	add	r0,r1,r3	; result in r3
        10'h085: pm_insn_o <= 16'h8025; // 	jmp	putc		; jump to putc to end it all
        10'h086: pm_insn_o <= 16'h419f; // 	set	#0x9f,r1	; 0x100 - 0x61 ('a')
        10'h087: pm_insn_o <= 16'h0101; // 	add	r0,r1,r1
        10'h088: pm_insn_o <= 16'h848d; // 	jmpc	convascii_gea	; Value is larger than or equal to 'a'
        10'h089: pm_insn_o <= 16'hffff; // 	nop
        10'h08a: pm_insn_o <= 16'h4007; // 	set	#0x7,r0		; ctrl g
        10'h08b: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h08c: pm_insn_o <= 16'h8077; // 	jmp	getnibble	; restart nibbleloop
        10'h08d: pm_insn_o <= 16'h4199; // 	set	#0x99,r1; 0x100 - 0x66 - 1 (0x66 = 'f')
        10'h08e: pm_insn_o <= 16'h0101; // 	add	r0,r1,r1
        10'h08f: pm_insn_o <= 16'h8494; // 	jmpc	invalidchar
        10'h090: pm_insn_o <= 16'hffff; // 	nop
        10'h091: pm_insn_o <= 16'h41a9; // 	set	#0xa9,r1	; -0x61+0xa
        10'h092: pm_insn_o <= 16'h0301; // 	add	r0,r1,r3	; result in r3
        10'h093: pm_insn_o <= 16'h8025; // 	jmp	putc
        10'h094: pm_insn_o <= 16'h4007; //  	set	#0x7,r0
        10'h095: pm_insn_o <= 16'h8625; //  	jsr	putc
        10'h096: pm_insn_o <= 16'h8077; // 	jmp	getnibble
        10'h097: pm_insn_o <= 16'h420f; // 	set	#0xf,r2 	; Mask out LSB nibble
        10'h098: pm_insn_o <= 16'h2202; // 	and	r0,r2,r2
        10'h099: pm_insn_o <= 16'h43f6; // 	set	#0xf6,r3
        10'h09a: pm_insn_o <= 16'h0323; // 	add	r2,r3,r3
        10'h09b: pm_insn_o <= 16'h84a0; // 	jmpc	convnibble_lsb_gtten ; Jump if r2 greater than 9
        10'h09c: pm_insn_o <= 16'hffff; // 	nop
        10'h09d: pm_insn_o <= 16'h4330; // 	set	#0x30,r3	; '0'
        10'h09e: pm_insn_o <= 16'h0123; // 	add	r2,r3,r1	; convert first nibble into '0'..'9'
        10'h09f: pm_insn_o <= 16'h80a2; // 	jmp	convnibble_msb
        10'h0a0: pm_insn_o <= 16'h4357; // 	set	#0x57,r3	; 'a'
        10'h0a1: pm_insn_o <= 16'h0123; // 	add	r2,r3,r1
        10'h0a2: pm_insn_o <= 16'h420f; // 	set	#0xf,r2		; mask out MSB nibble
        10'h0a3: pm_insn_o <= 16'h7000; // 	swap	r0,r0
        10'h0a4: pm_insn_o <= 16'h2202; // 	and	r0,r2,r2
        10'h0a5: pm_insn_o <= 16'h43f6; // 	set	#0xf6,r3
        10'h0a6: pm_insn_o <= 16'h0323; // 	add	r2,r3,r3
        10'h0a7: pm_insn_o <= 16'h84ac; // 	jmpc	convnibble_msb_gtten
        10'h0a8: pm_insn_o <= 16'hffff; // 	nop
        10'h0a9: pm_insn_o <= 16'h4330; // 	set	#0x30,r3	; '0'
        10'h0aa: pm_insn_o <= 16'h0023; // 	add	r2,r3,r0
        10'h0ab: pm_insn_o <= 16'h80ae; // 	jmp	convnibble_msb_done
        10'h0ac: pm_insn_o <= 16'h4357; // 	set	#0x57,r3	; 'a'
        10'h0ad: pm_insn_o <= 16'h0023; // 	add	r2,r3,r0
        10'h0ae: pm_insn_o <= 16'h3311; // 	or	r1,r1,r3	; move r1 to r3 FIXME - remove the need for this?
        10'h0af: pm_insn_o <= 16'h8800; // 	rts
        10'h0b0: pm_insn_o <= 16'h400d; // 	set	#0xd,r0
        10'h0b1: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h0b2: pm_insn_o <= 16'h400a; // 	set	#0xa,r0
        10'h0b3: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h0b4: pm_insn_o <= 16'h4001; // 	set	#0x1,r0
        10'h0b5: pm_insn_o <= 16'h0c0c; // 	add	r0,r12,r12
        10'h0b6: pm_insn_o <= 16'h0b0b; // 	add	r0,r11,r11
        10'h0b7: pm_insn_o <= 16'h84bb; // 	jmpc	nextrow_carry
        10'h0b8: pm_insn_o <= 16'hffff; // 	nop
        10'h0b9: pm_insn_o <= 16'h40ff; // 	set	#0xff,r0
        10'h0ba: pm_insn_o <= 16'h0c0c; // 	add	r0,r12,r12
        10'h0bb: pm_insn_o <= 16'h4508; // 	set	#0x8,r5
        10'h0bc: pm_insn_o <= 16'h4400; // 	set	#0x0,r4
        10'h0bd: pm_insn_o <= 16'h155c; // 	xor	r5,r12,r5
        10'h0be: pm_insn_o <= 16'h144b; // 	xor	r4,r11,r4
        10'h0bf: pm_insn_o <= 16'h3454; // 	or	r5,r4,r4
        10'h0c0: pm_insn_o <= 16'h820f; // 	jmpz	menuloop
        10'h0c1: pm_insn_o <= 16'hffff; // 	nop
        10'h0c2: pm_insn_o <= 16'h4d00; // 	set	LOW signalinfo,r13
        10'h0c3: pm_insn_o <= 16'h4700; // 	set	#0x0,r7
        10'h0c4: pm_insn_o <= 16'h4600; // 	set	#0x0,r6
        10'h0c5: pm_insn_o <= 16'h4500; // 	set	#0x0,r5
        10'h0c6: pm_insn_o <= 16'h4414; // 	set	#0x14,r4
        10'h0c7: pm_insn_o <= 16'h8730; // 	jsr	setwbaddr
        10'h0c8: pm_insn_o <= 16'h35cc; // 	or	r12,r12,r5
        10'h0c9: pm_insn_o <= 16'h34bb; // 	or	r11,r11,r4
        10'h0ca: pm_insn_o <= 16'h8732; // 	jsr	setwbdata
        10'h0cb: pm_insn_o <= 16'h872b; // 	jsr	write_to_wb
        10'h0cc: pm_insn_o <= 16'h80d3; // 	jmp	handle_logicanalyzer_mainloop
        10'h0cd: pm_insn_o <= 16'h4300; // 	set	LOW signalnames,r3
        10'h0ce: pm_insn_o <= 16'h4406; // 	set	HIGH signalnames,r4
        10'h0cf: pm_insn_o <= 16'h87d3; // 	jsr	puts
        10'h0d0: pm_insn_o <= 16'h4b00; // 	set	#0x0,r11
        10'h0d1: pm_insn_o <= 16'h4c00; // 	set	#0x0,r12	;  Entry to display...
        10'h0d2: pm_insn_o <= 16'h80c2; // 	jmp	nextrow_setup
        10'h0d3: pm_insn_o <= 16'h4009; // 	set	#0x9,r0		; tab
        10'h0d4: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h0d5: pm_insn_o <= 16'h4104; // 	set	HIGH signalinfo,r1
        10'h0d6: pm_insn_o <= 16'h6e1d; // 	ld	r1,r13,r14
        10'h0d7: pm_insn_o <= 16'h6e1d; // 	ld	r1,r13,r14
        10'h0d8: pm_insn_o <= 16'h4001; // 	set	#0x1,r0
        10'h0d9: pm_insn_o <= 16'h0d0d; // 	add	r0,r13,r13
        10'h0da: pm_insn_o <= 16'h6f1d; // 	ld	r1,r13,r15
        10'h0db: pm_insn_o <= 16'h6f1d; // 	ld	r1,r13,r15
        10'h0dc: pm_insn_o <= 16'h0d0d; // 	add	r0,r13,r13
        10'h0dd: pm_insn_o <= 16'h3eee; // 	or	r14,r14,r14
        10'h0de: pm_insn_o <= 16'h82b0; // 	jmpz	logicanalyzer_nextrow	; Finished (well, not really...)
        10'h0df: pm_insn_o <= 16'hffff; // 	nop
        10'h0e0: pm_insn_o <= 16'h4900; // 	set	#0x0,r9
        10'h0e1: pm_insn_o <= 16'h38ff; // 	or	r15,r15,r8
        10'h0e2: pm_insn_o <= 16'h8702; // 	jsr	getbit_from_analyzer
        10'h0e3: pm_insn_o <= 16'h0999; // 	add	r9,r9,r9
        10'h0e4: pm_insn_o <= 16'h3989; // 	or	r8,r9,r9
        10'h0e5: pm_insn_o <= 16'h40ff; // 	set	#0xff,r0
        10'h0e6: pm_insn_o <= 16'h0f0f; // 	add	r0,r15,r15
        10'h0e7: pm_insn_o <= 16'h0e0e; // 	add	r0,r14,r14
        10'h0e8: pm_insn_o <= 16'h4003; // 	set	#0x3,r0
        10'h0e9: pm_insn_o <= 16'h200e; // 	and	r0,r14,r0
        10'h0ea: pm_insn_o <= 16'h82f0; // 	jmpz	logicloop_printnibble
        10'h0eb: pm_insn_o <= 16'hffff; // 	nop
        10'h0ec: pm_insn_o <= 16'h3eee; // 	or	r14,r14,r14
        10'h0ed: pm_insn_o <= 16'h82d3; // 	jmpz	handle_logicanalyzer_mainloop
        10'h0ee: pm_insn_o <= 16'hffff; // 	nop
        10'h0ef: pm_insn_o <= 16'h80e1; // 	jmp	logicloop
        10'h0f0: pm_insn_o <= 16'h3099; // 	or	r9,r9,r0
        10'h0f1: pm_insn_o <= 16'h8697; // 	jsr	convnibble
        10'h0f2: pm_insn_o <= 16'h3033; // 	or	r3,r3,r0
        10'h0f3: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h0f4: pm_insn_o <= 16'h4900; // 	set	#0x0,r9
        10'h0f5: pm_insn_o <= 16'h80ec; // 	jmp	logicloop_continue
        10'h0f6: pm_insn_o <= 16'h4018; // 	set	#0x18,r0
        10'h0f7: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h0f8: pm_insn_o <= 16'h45f1; // 	set	#0xf1,r5	; Read, sel is 0xf
        10'h0f9: pm_insn_o <= 16'h9150; // 	out1	r5
        10'h0fa: pm_insn_o <= 16'h8800; // 	rts
        10'h0fb: pm_insn_o <= 16'h4101; // 	set	#0x1,r1
        10'h0fc: pm_insn_o <= 16'h0000; // 	add	r0,r0,r0
        10'h0fd: pm_insn_o <= 16'h8500; // 	jmpc	rol1_carry
        10'h0fe: pm_insn_o <= 16'hffff; // 	nop
        10'h0ff: pm_insn_o <= 16'h8800; // 	rts
        10'h100: pm_insn_o <= 16'h0001; // 	add	r0,r1,r0
        10'h101: pm_insn_o <= 16'h8800; // 	rts
        10'h102: pm_insn_o <= 16'h41e0; // 	set	#0xe0,r1
        10'h103: pm_insn_o <= 16'h2081; // 	and	r8,r1,r0	; r0 contains the address to read from logicanalyzer
        10'h104: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h105: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h106: pm_insn_o <= 16'h86fb; // 	jsr	rol1		
        10'h107: pm_insn_o <= 16'h0000; // 	add	r0,r0,r0	; Multiply it with 2
        10'h108: pm_insn_o <= 16'h0000; // 	add	r0,r0,r0
        10'h109: pm_insn_o <= 16'h4140; // 	set	#0x40,r1
        10'h10a: pm_insn_o <= 16'h0401; // 	add	r0,r1,r4	; Add the offset to logic analyzer port (0x40) to it
        10'h10b: pm_insn_o <= 16'h4500; // 	set	#0x0,r5
        10'h10c: pm_insn_o <= 16'h4600; // 	set	#0x0,r6
        10'h10d: pm_insn_o <= 16'h4700; // 	set	#0x0,r7
        10'h10e: pm_insn_o <= 16'h4010; // 	set	#0x10,r0	; Set wishbone address 
        10'h10f: pm_insn_o <= 16'h8655; // 	jsr	setport		; r4-r7 -> port 0x10 => wb addr
        10'h110: pm_insn_o <= 16'h86f6; // 	jsr	wishbone_do_read
        10'h111: pm_insn_o <= 16'h4118; // 	set	#0x18,r1	; Byte to read
        10'h112: pm_insn_o <= 16'h2081; // 	and	r8,r1,r0	
        10'h113: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h114: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h115: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h116: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h117: pm_insn_o <= 16'h86fb; // 	jsr	rol1		; r0 now contains the byte to read from logicanalyzer
        10'h118: pm_insn_o <= 16'h4114; // 	set	#0x14,r1	; offset to WB master peripheral
        10'h119: pm_insn_o <= 16'h0101; // 	add	r0,r1,r1
        10'h11a: pm_insn_o <= 16'h9010; // 	out0	r1
        10'h11b: pm_insn_o <= 16'h4107; // 	set	#0x7,r1
        10'h11c: pm_insn_o <= 16'h2081; // 	and	r8,r1,r0	; r0 contains the bitnumber we are interested in
        10'h11d: pm_insn_o <= 16'h5800; // 	in2	r8		; r8 now contains the byte we are interested in
        10'h11e: pm_insn_o <= 16'h43ff; // 	set	#0xff,r3
        10'h11f: pm_insn_o <= 16'h4201; // 	set	#0x1,r2		; mask
        10'h120: pm_insn_o <= 16'h3000; // 	or	r0,r0,r0
        10'h121: pm_insn_o <= 16'h8326; // 	jmpz	getbit_loopend
        10'h122: pm_insn_o <= 16'hffff; // 	nop
        10'h123: pm_insn_o <= 16'h0003; // 	add	r0,r3,r0	; r0--
        10'h124: pm_insn_o <= 16'h0222; // 	add	r2,r2,r2	; r2 = r2 << 1
        10'h125: pm_insn_o <= 16'h8120; // 	jmp	getbit_loopstart
        10'h126: pm_insn_o <= 16'h2828; // 	and	r2,r8,r8	; r8 is now masked
        10'h127: pm_insn_o <= 16'h832a; // 	jmpz	getbit_iszero
        10'h128: pm_insn_o <= 16'hffff; // 	nop
        10'h129: pm_insn_o <= 16'h4801; // 	set	#0x1,r8
        10'h12a: pm_insn_o <= 16'h8800; // 	rts
        10'h12b: pm_insn_o <= 16'h4018; // 	set	#0x18,r0
        10'h12c: pm_insn_o <= 16'h41f9; // 	set	#0xf9,r1
        10'h12d: pm_insn_o <= 16'h9000; // 	out0	r0
        10'h12e: pm_insn_o <= 16'h9110; // 	out1	r1
        10'h12f: pm_insn_o <= 16'h8800; // 	rts
        10'h130: pm_insn_o <= 16'h4010; // 	set	#0x10,r0
        10'h131: pm_insn_o <= 16'h8055; // 	jmp	setport
        10'h132: pm_insn_o <= 16'h4014; // 	set	#0x14,r0
        10'h133: pm_insn_o <= 16'h8055; // 	jmp	setport
        10'h134: pm_insn_o <= 16'h4700; // 	set	#0x0,r7
        10'h135: pm_insn_o <= 16'h4600; // 	set	#0x0,r6
        10'h136: pm_insn_o <= 16'h4500; // 	set	#0x0,r5
        10'h137: pm_insn_o <= 16'h4420; // 	set	#0x20,r4
        10'h138: pm_insn_o <= 16'h8730; // 	jsr	setwbaddr
        10'h139: pm_insn_o <= 16'h4400; // 	set	#0x0,r4
        10'h13a: pm_insn_o <= 16'h8732; // 	jsr	setwbdata
        10'h13b: pm_insn_o <= 16'h872b; // 	jsr	write_to_wb	;  Stop tracer machine
        10'h13c: pm_insn_o <= 16'h4700; // 	set	#0x0,r7
        10'h13d: pm_insn_o <= 16'h4600; // 	set	#0x0,r6
        10'h13e: pm_insn_o <= 16'h4500; // 	set	#0x0,r5
        10'h13f: pm_insn_o <= 16'h4400; // 	set	#0x0,r4
        10'h140: pm_insn_o <= 16'h8730; // 	jsr	setwbaddr
        10'h141: pm_insn_o <= 16'h4401; // 	set	#0x1,r4
        10'h142: pm_insn_o <= 16'h8732; // 	jsr	setwbdata
        10'h143: pm_insn_o <= 16'h872b; // 	jsr	write_to_wb
        10'h144: pm_insn_o <= 16'h86f6; // 	jsr	wishbone_do_read
        10'h145: pm_insn_o <= 16'h4014; // 	set	#0x14,r0
        10'h146: pm_insn_o <= 16'h8662; // 	jsr	getport
        10'h147: pm_insn_o <= 16'h3444; // 	or	r4,r4,r4
        10'h148: pm_insn_o <= 16'h8344; // 	jmpz	handle_trigger_wait
        10'h149: pm_insn_o <= 16'h4330; // 	set	LOW triggermessage,r3
        10'h14a: pm_insn_o <= 16'h4405; // 	set	HIGH triggermessage,r4
        10'h14b: pm_insn_o <= 16'h800e; // 	jmp	greetloop
        10'h14c: pm_insn_o <= 16'h4201; // 	set	#0x1,r2
        10'h14d: pm_insn_o <= 16'h43ff; // 	set	#0xff,r3
        10'h14e: pm_insn_o <= 16'h3000; // 	or	r0,r0,r0
        10'h14f: pm_insn_o <= 16'h8354; // 	jmpz	createbitmask_end
        10'h150: pm_insn_o <= 16'hffff; // 	nop
        10'h151: pm_insn_o <= 16'h0003; // 	add	r0,r3,r0	; r0--
        10'h152: pm_insn_o <= 16'h0222; // 	add	r2,r2,r2	; r2 = r2 << 1
        10'h153: pm_insn_o <= 16'h814e; // 	jmp	createbitmask_loop
        10'h154: pm_insn_o <= 16'h8800; // 	rts
        10'h155: pm_insn_o <= 16'h4700; // 	set	#0x00,r7
        10'h156: pm_insn_o <= 16'h4600; // 	set	#0x00,r6
        10'h157: pm_insn_o <= 16'h4500; // 	set	#0x00,r5
        10'h158: pm_insn_o <= 16'h34bb; // 	or	r11,r11,r4
        10'h159: pm_insn_o <= 16'h41e0; // 	set	#0xe0,r1
        10'h15a: pm_insn_o <= 16'h2081; // 	and	r8,r1,r0
        10'h15b: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h15c: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h15d: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h15e: pm_insn_o <= 16'h0000; // 	add	r0,r0,r0
        10'h15f: pm_insn_o <= 16'h0000; // 	add	r0,r0,r0
        10'h160: pm_insn_o <= 16'h0404; // 	add	r0,r4,r4	; r7-r4 now contains WB word for matchbit
        10'h161: pm_insn_o <= 16'h8730; // 	jsr	setwbaddr
        10'h162: pm_insn_o <= 16'h86f6; // 	jsr	wishbone_do_read
        10'h163: pm_insn_o <= 16'h4118; // 	set	#0x18,r1	; Byte to read
        10'h164: pm_insn_o <= 16'h2081; // 	and	r8,r1,r0	
        10'h165: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h166: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h167: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h168: pm_insn_o <= 16'h86fb; // 	jsr	rol1
        10'h169: pm_insn_o <= 16'h86fb; // 	jsr	rol1		; r0 now contains the byte to read from logicanalyzer
        10'h16a: pm_insn_o <= 16'h4114; // 	set	#0x14,r1	; offset to WB master peripheral
        10'h16b: pm_insn_o <= 16'h0a01; // 	add	r0,r1,r10	; Save port offset in r10
        10'h16c: pm_insn_o <= 16'h90a0; // 	out0	r10
        10'h16d: pm_insn_o <= 16'h5400; // 	in2	r4		; r4 contains the byte we want to mask
        10'h16e: pm_insn_o <= 16'h4107; // 	set	#0x7,r1
        10'h16f: pm_insn_o <= 16'h2081; // 	and	r8,r1,r0	; r0 contains the bitnumber we are interested in
        10'h170: pm_insn_o <= 16'h874c; // 	jsr	createbitmask
        10'h171: pm_insn_o <= 16'h43ff; // 	set	#0xff,r3
        10'h172: pm_insn_o <= 16'h1323; // 	xor	r2,r3,r3	; r3 now contains inverted mask for anding
        10'h173: pm_insn_o <= 16'h2443; // 	and	r4,r3,r4	; r4 is now cleared
        10'h174: pm_insn_o <= 16'h3999; // 	or	r9,r9,r9	; set flags
        10'h175: pm_insn_o <= 16'h8378; // 	jmpz	setbit_writeback
        10'h176: pm_insn_o <= 16'hffff; // 	nop
        10'h177: pm_insn_o <= 16'h3442; // 	or	r4,r2,r4	; r9 now contains correct byte value
        10'h178: pm_insn_o <= 16'h3944; // 	or	r4,r4,r9	; Save byte in r9
        10'h179: pm_insn_o <= 16'h4014; // 	set	#0x14,r0
        10'h17a: pm_insn_o <= 16'h8662; // 	jsr	getport		; Read port data
        10'h17b: pm_insn_o <= 16'h4014; // 	set	#0x14,r0
        10'h17c: pm_insn_o <= 16'h8655; // 	jsr	setport		; Write it back
        10'h17d: pm_insn_o <= 16'h90a0; // 	out0	r10		; Update this particular byte
        10'h17e: pm_insn_o <= 16'h9190; // 	out1	r9
        10'h17f: pm_insn_o <= 16'h812b; // 	jmp	write_to_wb
        10'h180: pm_insn_o <= 16'h4300; // 	set	LOW signalnames,r3
        10'h181: pm_insn_o <= 16'h4406; // 	set	HIGH signalnames,r4
        10'h182: pm_insn_o <= 16'h87d3; // 	jsr	puts
        10'h183: pm_insn_o <= 16'h4b00; // 	set	#0x0,r11
        10'h184: pm_insn_o <= 16'h4000; // 	set	#0x0,r0
        10'h185: pm_insn_o <= 16'h10b0; // 	xor	r11,r0,r0
        10'h186: pm_insn_o <= 16'h8390; // 	jmpz	handle_settrigger_setval
        10'h187: pm_insn_o <= 16'h400c; // 	set	#0xc,r0
        10'h188: pm_insn_o <= 16'h10b0; // 	xor	r11,r0,r0
        10'h189: pm_insn_o <= 16'h838b; // 	jmpz	handle_settrigger_setmask
        10'h18a: pm_insn_o <= 16'h800f; // 	jmp	menuloop	; Exit handle_settrigger
        10'h18b: pm_insn_o <= 16'h4b04; // 	set	#0x4,r11
        10'h18c: pm_insn_o <= 16'h4322; // 	set	LOW maskvalstring,r3
        10'h18d: pm_insn_o <= 16'h4405; // 	set	HIGH maskvalstring,r4
        10'h18e: pm_insn_o <= 16'h87d3; // 	jsr	puts
        10'h18f: pm_insn_o <= 16'h8194; // 	jmp	handle_settrigger_main
        10'h190: pm_insn_o <= 16'h4314; // 	set	LOW trigvalstring,r3
        10'h191: pm_insn_o <= 16'h4405; // 	set	HIGH trigvalstring,r4
        10'h192: pm_insn_o <= 16'h87d3; // 	jsr	puts
        10'h193: pm_insn_o <= 16'h4b0c; // 	set	#0xc,r11
        10'h194: pm_insn_o <= 16'h4d00; // 	set	LOW signalinfo,r13 ;r13 contains pointer to current
        10'h195: pm_insn_o <= 16'h4009; // 	set	#0x9,r0		; '\t'
        10'h196: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h197: pm_insn_o <= 16'h4104; // 	set	HIGH signalinfo,r1
        10'h198: pm_insn_o <= 16'h6e1d; // 	ld	r1,r13,r14	   
        10'h199: pm_insn_o <= 16'h6e1d; // 	ld	r1,r13,r14	   ;r14 contains length of current entry
        10'h19a: pm_insn_o <= 16'h3eee; // 	or	r14,r14,r14
        10'h19b: pm_insn_o <= 16'h8384; // 	jmpz	handle_settrigger_setvalormask	; No more entry
        10'h19c: pm_insn_o <= 16'hffff; // 	nop
        10'h19d: pm_insn_o <= 16'h4001; // 	set	#0x1,r0
        10'h19e: pm_insn_o <= 16'h0d0d; // 	add	r0,r13,r13
        10'h19f: pm_insn_o <= 16'h6f1d; // 	ld	r1,r13,r15	
        10'h1a0: pm_insn_o <= 16'h6f1d; // 	ld	r1,r13,r15	; r15 contains bit offset of current entry
        10'h1a1: pm_insn_o <= 16'h0d0d; // 	add	r0,r13,r13	; r13 points to next entry
        10'h1a2: pm_insn_o <= 16'h3eee; // 	or	r14,r14,r14
        10'h1a3: pm_insn_o <= 16'h8395; // 	jmpz	handle_settrigger_nextentry	; No more entry
        10'h1a4: pm_insn_o <= 16'hffff; // 	nop
        10'h1a5: pm_insn_o <= 16'h8677; // 	jsr	getnibble	; r3 contains input
        10'h1a6: pm_insn_o <= 16'h3c33; // 	or	r3,r3,r12
        10'h1a7: pm_insn_o <= 16'h4203; // 	set	#0x3,r2
        10'h1a8: pm_insn_o <= 16'h222e; // 	and	r2,r14,r2	; r2 contains length & 3
        10'h1a9: pm_insn_o <= 16'h4900; // 	set	#0x0,r9
        10'h1aa: pm_insn_o <= 16'h1992; // 	xor	r9,r2,r9	; (length & 3) == 0 ?
        10'h1ab: pm_insn_o <= 16'h83b5; // 	jmpz	handle_settrigger_use4
        10'h1ac: pm_insn_o <= 16'h4903; // 	set	#0x3,r9
        10'h1ad: pm_insn_o <= 16'h1992; // 	xor	r9,r2,r9	; (length & 3) == 3 ?
        10'h1ae: pm_insn_o <= 16'h83bc; // 	jmpz	handle_settrigger_use3
        10'h1af: pm_insn_o <= 16'h4902; // 	set	#0x2,r9
        10'h1b0: pm_insn_o <= 16'h1992; // 	xor	r9,r2,r9	; (length & 3) == 2 ?
        10'h1b1: pm_insn_o <= 16'h83c3; // 	jmpz	handle_settrigger_use2
        10'h1b2: pm_insn_o <= 16'h4901; // 	set	#0x1,r9
        10'h1b3: pm_insn_o <= 16'h1992; // 	xor	r9,r2,r9	; (length & 3) == 1 ?
        10'h1b4: pm_insn_o <= 16'h83ca; // 	jmpz	handle_settrigger_use1
        10'h1b5: pm_insn_o <= 16'h4008; // 	set	#0x8,r0
        10'h1b6: pm_insn_o <= 16'h290c; // 	and	r0,r12,r9
        10'h1b7: pm_insn_o <= 16'h38ff; // 	or	r15,r15,r8
        10'h1b8: pm_insn_o <= 16'h8755; // 	jsr	setbit
        10'h1b9: pm_insn_o <= 16'h4aff; // 	set	#0xff,r10	; r10 = -1
        10'h1ba: pm_insn_o <= 16'h0eea; // 	add	r14,r10,r14
        10'h1bb: pm_insn_o <= 16'h0ffa; // 	add	r15,r10,r15
        10'h1bc: pm_insn_o <= 16'h4004; // 	set	#0x4,r0
        10'h1bd: pm_insn_o <= 16'h290c; // 	and	r0,r12,r9
        10'h1be: pm_insn_o <= 16'h38ff; // 	or	r15,r15,r8
        10'h1bf: pm_insn_o <= 16'h8755; // 	jsr	setbit
        10'h1c0: pm_insn_o <= 16'h4aff; // 	set	#0xff,r10	; r10 = -1
        10'h1c1: pm_insn_o <= 16'h0eea; // 	add	r14,r10,r14
        10'h1c2: pm_insn_o <= 16'h0ffa; // 	add	r15,r10,r15
        10'h1c3: pm_insn_o <= 16'h4002; // 	set	#0x2,r0
        10'h1c4: pm_insn_o <= 16'h290c; // 	and	r0,r12,r9
        10'h1c5: pm_insn_o <= 16'h38ff; // 	or	r15,r15,r8
        10'h1c6: pm_insn_o <= 16'h8755; // 	jsr	setbit
        10'h1c7: pm_insn_o <= 16'h4aff; // 	set	#0xff,r10	; r10 = -1
        10'h1c8: pm_insn_o <= 16'h0eea; // 	add	r14,r10,r14
        10'h1c9: pm_insn_o <= 16'h0ffa; // 	add	r15,r10,r15
        10'h1ca: pm_insn_o <= 16'h4001; // 	set	#0x1,r0
        10'h1cb: pm_insn_o <= 16'h290c; // 	and	r0,r12,r9
        10'h1cc: pm_insn_o <= 16'h38ff; // 	or	r15,r15,r8
        10'h1cd: pm_insn_o <= 16'h8755; // 	jsr	setbit
        10'h1ce: pm_insn_o <= 16'h4aff; // 	set	#0xff,r10	; r10 = -1
        10'h1cf: pm_insn_o <= 16'h0eea; // 	add	r14,r10,r14
        10'h1d0: pm_insn_o <= 16'h0ffa; // 	add	r15,r10,r15
        10'h1d1: pm_insn_o <= 16'h81a2; // 	jmp	handle_settrigger_nextnibble
        10'h1d2: pm_insn_o <= 16'h800f; // 	jmp	menuloop
        10'h1d3: pm_insn_o <= 16'h6043; // 	ld	r4,r3,r0
        10'h1d4: pm_insn_o <= 16'h6043; // 	ld	r4,r3,r0
        10'h1d5: pm_insn_o <= 16'h3000; // 	or	r0,r0,r0
        10'h1d6: pm_insn_o <= 16'h83dc; // 	jmpz	end_puts
        10'h1d7: pm_insn_o <= 16'hffff; // 	nop
        10'h1d8: pm_insn_o <= 16'h8625; // 	jsr	putc
        10'h1d9: pm_insn_o <= 16'h4001; // 	set	#0x01,r0
        10'h1da: pm_insn_o <= 16'h0303; // 	add	r0,r3,r3	;charptr++
        10'h1db: pm_insn_o <= 16'h81d3; // 	jmp	puts
        10'h1dc: pm_insn_o <= 16'h8800; // 	rts
        10'h1dd: pm_insn_o <= 16'h0000;
        10'h1de: pm_insn_o <= 16'h0000;
        10'h1df: pm_insn_o <= 16'h0000;
        10'h1e0: pm_insn_o <= 16'h0000;
        10'h1e1: pm_insn_o <= 16'h0000;
        10'h1e2: pm_insn_o <= 16'h0000;
        10'h1e3: pm_insn_o <= 16'h0000;
        10'h1e4: pm_insn_o <= 16'h0000;
        10'h1e5: pm_insn_o <= 16'h0000;
        10'h1e6: pm_insn_o <= 16'h0000;
        10'h1e7: pm_insn_o <= 16'h0000;
        10'h1e8: pm_insn_o <= 16'h0000;
        10'h1e9: pm_insn_o <= 16'h0000;
        10'h1ea: pm_insn_o <= 16'h0000;
        10'h1eb: pm_insn_o <= 16'h0000;
        10'h1ec: pm_insn_o <= 16'h0000;
        10'h1ed: pm_insn_o <= 16'h0000;
        10'h1ee: pm_insn_o <= 16'h0000;
        10'h1ef: pm_insn_o <= 16'h0000;
        10'h1f0: pm_insn_o <= 16'h0000;
        10'h1f1: pm_insn_o <= 16'h0000;
        10'h1f2: pm_insn_o <= 16'h0000;
        10'h1f3: pm_insn_o <= 16'h0000;
        10'h1f4: pm_insn_o <= 16'h0000;
        10'h1f5: pm_insn_o <= 16'h0000;
        10'h1f6: pm_insn_o <= 16'h0000;
        10'h1f7: pm_insn_o <= 16'h0000;
        10'h1f8: pm_insn_o <= 16'h0000;
        10'h1f9: pm_insn_o <= 16'h0000;
        10'h1fa: pm_insn_o <= 16'h0000;
        10'h1fb: pm_insn_o <= 16'h0000;
        10'h1fc: pm_insn_o <= 16'h0000;
        10'h1fd: pm_insn_o <= 16'h0000;
        10'h1fe: pm_insn_o <= 16'h0000;
        10'h1ff: pm_insn_o <= 16'h0000;
        10'h200: pm_insn_o <= 16'h070e; // 	dw	0x070e
        10'h201: pm_insn_o <= 16'h0807; // 	dw	0x0807
        10'h202: pm_insn_o <= 16'h0000; // 	dw	0x0000
        10'h203: pm_insn_o <= 16'h0000; // 	dw	0x0000
        10'h204: pm_insn_o <= 16'h0000;
        10'h205: pm_insn_o <= 16'h0000;
        10'h206: pm_insn_o <= 16'h0000;
        10'h207: pm_insn_o <= 16'h0000;
        10'h208: pm_insn_o <= 16'h0000;
        10'h209: pm_insn_o <= 16'h0000;
        10'h20a: pm_insn_o <= 16'h0000;
        10'h20b: pm_insn_o <= 16'h0000;
        10'h20c: pm_insn_o <= 16'h0000;
        10'h20d: pm_insn_o <= 16'h0000;
        10'h20e: pm_insn_o <= 16'h0000;
        10'h20f: pm_insn_o <= 16'h0000;
        10'h210: pm_insn_o <= 16'h0000;
        10'h211: pm_insn_o <= 16'h0000;
        10'h212: pm_insn_o <= 16'h0000;
        10'h213: pm_insn_o <= 16'h0000;
        10'h214: pm_insn_o <= 16'h0000;
        10'h215: pm_insn_o <= 16'h0000;
        10'h216: pm_insn_o <= 16'h0000;
        10'h217: pm_insn_o <= 16'h0000;
        10'h218: pm_insn_o <= 16'h0000;
        10'h219: pm_insn_o <= 16'h0000;
        10'h21a: pm_insn_o <= 16'h0000;
        10'h21b: pm_insn_o <= 16'h0000;
        10'h21c: pm_insn_o <= 16'h0000;
        10'h21d: pm_insn_o <= 16'h0000;
        10'h21e: pm_insn_o <= 16'h0000;
        10'h21f: pm_insn_o <= 16'h0000;
        10'h220: pm_insn_o <= 16'h0000;
        10'h221: pm_insn_o <= 16'h0000;
        10'h222: pm_insn_o <= 16'h0000;
        10'h223: pm_insn_o <= 16'h0000;
        10'h224: pm_insn_o <= 16'h0000;
        10'h225: pm_insn_o <= 16'h0000;
        10'h226: pm_insn_o <= 16'h0000;
        10'h227: pm_insn_o <= 16'h0000;
        10'h228: pm_insn_o <= 16'h0000;
        10'h229: pm_insn_o <= 16'h0000;
        10'h22a: pm_insn_o <= 16'h0000;
        10'h22b: pm_insn_o <= 16'h0000;
        10'h22c: pm_insn_o <= 16'h0000;
        10'h22d: pm_insn_o <= 16'h0000;
        10'h22e: pm_insn_o <= 16'h0000;
        10'h22f: pm_insn_o <= 16'h0000;
        10'h230: pm_insn_o <= 16'h0000;
        10'h231: pm_insn_o <= 16'h0000;
        10'h232: pm_insn_o <= 16'h0000;
        10'h233: pm_insn_o <= 16'h0000;
        10'h234: pm_insn_o <= 16'h0000;
        10'h235: pm_insn_o <= 16'h0000;
        10'h236: pm_insn_o <= 16'h0000;
        10'h237: pm_insn_o <= 16'h0000;
        10'h238: pm_insn_o <= 16'h0000;
        10'h239: pm_insn_o <= 16'h0000;
        10'h23a: pm_insn_o <= 16'h0000;
        10'h23b: pm_insn_o <= 16'h0000;
        10'h23c: pm_insn_o <= 16'h0000;
        10'h23d: pm_insn_o <= 16'h0000;
        10'h23e: pm_insn_o <= 16'h0000;
        10'h23f: pm_insn_o <= 16'h0000;
        10'h240: pm_insn_o <= 16'h0000;
        10'h241: pm_insn_o <= 16'h0000;
        10'h242: pm_insn_o <= 16'h0000;
        10'h243: pm_insn_o <= 16'h0000;
        10'h244: pm_insn_o <= 16'h0000;
        10'h245: pm_insn_o <= 16'h0000;
        10'h246: pm_insn_o <= 16'h0000;
        10'h247: pm_insn_o <= 16'h0000;
        10'h248: pm_insn_o <= 16'h0000;
        10'h249: pm_insn_o <= 16'h0000;
        10'h24a: pm_insn_o <= 16'h0000;
        10'h24b: pm_insn_o <= 16'h0000;
        10'h24c: pm_insn_o <= 16'h0000;
        10'h24d: pm_insn_o <= 16'h0000;
        10'h24e: pm_insn_o <= 16'h0000;
        10'h24f: pm_insn_o <= 16'h0000;
        10'h250: pm_insn_o <= 16'h0000;
        10'h251: pm_insn_o <= 16'h0000;
        10'h252: pm_insn_o <= 16'h0000;
        10'h253: pm_insn_o <= 16'h0000;
        10'h254: pm_insn_o <= 16'h0000;
        10'h255: pm_insn_o <= 16'h0000;
        10'h256: pm_insn_o <= 16'h0000;
        10'h257: pm_insn_o <= 16'h0000;
        10'h258: pm_insn_o <= 16'h0000;
        10'h259: pm_insn_o <= 16'h0000;
        10'h25a: pm_insn_o <= 16'h0000;
        10'h25b: pm_insn_o <= 16'h0000;
        10'h25c: pm_insn_o <= 16'h0000;
        10'h25d: pm_insn_o <= 16'h0000;
        10'h25e: pm_insn_o <= 16'h0000;
        10'h25f: pm_insn_o <= 16'h0000;
        10'h260: pm_insn_o <= 16'h0000;
        10'h261: pm_insn_o <= 16'h0000;
        10'h262: pm_insn_o <= 16'h0000;
        10'h263: pm_insn_o <= 16'h0000;
        10'h264: pm_insn_o <= 16'h0000;
        10'h265: pm_insn_o <= 16'h0000;
        10'h266: pm_insn_o <= 16'h0000;
        10'h267: pm_insn_o <= 16'h0000;
        10'h268: pm_insn_o <= 16'h0000;
        10'h269: pm_insn_o <= 16'h0000;
        10'h26a: pm_insn_o <= 16'h0000;
        10'h26b: pm_insn_o <= 16'h0000;
        10'h26c: pm_insn_o <= 16'h0000;
        10'h26d: pm_insn_o <= 16'h0000;
        10'h26e: pm_insn_o <= 16'h0000;
        10'h26f: pm_insn_o <= 16'h0000;
        10'h270: pm_insn_o <= 16'h0000;
        10'h271: pm_insn_o <= 16'h0000;
        10'h272: pm_insn_o <= 16'h0000;
        10'h273: pm_insn_o <= 16'h0000;
        10'h274: pm_insn_o <= 16'h0000;
        10'h275: pm_insn_o <= 16'h0000;
        10'h276: pm_insn_o <= 16'h0000;
        10'h277: pm_insn_o <= 16'h0000;
        10'h278: pm_insn_o <= 16'h0000;
        10'h279: pm_insn_o <= 16'h0000;
        10'h27a: pm_insn_o <= 16'h0000;
        10'h27b: pm_insn_o <= 16'h0000;
        10'h27c: pm_insn_o <= 16'h0000;
        10'h27d: pm_insn_o <= 16'h0000;
        10'h27e: pm_insn_o <= 16'h0000;
        10'h27f: pm_insn_o <= 16'h0000;
        10'h280: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a		; \r\n
        10'h281: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a		; \r\n
        10'h282: pm_insn_o <= 16'h2a2a; // 	dw	0x2a2a		; **
        10'h283: pm_insn_o <= 16'h2a20; // 	dw	0x2a20		; *
        10'h284: pm_insn_o <= 16'h4145; // 	dw	0x4145		; AE
        10'h285: pm_insn_o <= 16'h2044; // 	dw	0x2044		;  D
        10'h286: pm_insn_o <= 16'h6562; // 	dw	0x6562		; eb
        10'h287: pm_insn_o <= 16'h7567; // 	dw	0x7567		; ug
        10'h288: pm_insn_o <= 16'h2049; // 	dw	0x2049		;  I
        10'h289: pm_insn_o <= 16'h4600; // 	dw	0x4600		; F\0
        10'h28a: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a		; \r\n
        10'h28b: pm_insn_o <= 16'h5472; // 	dw	0x5472		;
        10'h28c: pm_insn_o <= 16'h6967; // 	dw	0x6967
        10'h28d: pm_insn_o <= 16'h7661; // 	dw	0x7661
        10'h28e: pm_insn_o <= 16'h6c3a; // 	dw	0x6c3a
        10'h28f: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a		; \r\n
        10'h290: pm_insn_o <= 16'h0000; // 	dw	0x0000
        10'h291: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a		; \r\n
        10'h292: pm_insn_o <= 16'h4d61; // 	dw	0x4d61
        10'h293: pm_insn_o <= 16'h736b; // 	dw	0x736b
        10'h294: pm_insn_o <= 16'h7661; // 	dw	0x7661
        10'h295: pm_insn_o <= 16'h6c3a; // 	dw	0x6c3a
        10'h296: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a		; \r\n
        10'h297: pm_insn_o <= 16'h0000; // 	dw	0x0000
        10'h298: pm_insn_o <= 16'h5761; // 	dw	0x5761
        10'h299: pm_insn_o <= 16'h6974; // 	dw	0x6974
        10'h29a: pm_insn_o <= 16'h696e; // 	dw	0x696e
        10'h29b: pm_insn_o <= 16'h6720; // 	dw	0x6720
        10'h29c: pm_insn_o <= 16'h666f; // 	dw	0x666f
        10'h29d: pm_insn_o <= 16'h7220; // 	dw	0x7220
        10'h29e: pm_insn_o <= 16'h7472; // 	dw	0x7472
        10'h29f: pm_insn_o <= 16'h6967; // 	dw	0x6967
        10'h2a0: pm_insn_o <= 16'h6765; // 	dw	0x6765
        10'h2a1: pm_insn_o <= 16'h722e; // 	dw	0x722e
        10'h2a2: pm_insn_o <= 16'h2e2e; // 	dw	0x2e2e
        10'h2a3: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a
        10'h2a4: pm_insn_o <= 16'h0000; // 	dw	0x0000
        10'h2a5: pm_insn_o <= 16'h0000;
        10'h2a6: pm_insn_o <= 16'h0000;
        10'h2a7: pm_insn_o <= 16'h0000;
        10'h2a8: pm_insn_o <= 16'h0000;
        10'h2a9: pm_insn_o <= 16'h0000;
        10'h2aa: pm_insn_o <= 16'h0000;
        10'h2ab: pm_insn_o <= 16'h0000;
        10'h2ac: pm_insn_o <= 16'h0000;
        10'h2ad: pm_insn_o <= 16'h0000;
        10'h2ae: pm_insn_o <= 16'h0000;
        10'h2af: pm_insn_o <= 16'h0000;
        10'h2b0: pm_insn_o <= 16'h0000;
        10'h2b1: pm_insn_o <= 16'h0000;
        10'h2b2: pm_insn_o <= 16'h0000;
        10'h2b3: pm_insn_o <= 16'h0000;
        10'h2b4: pm_insn_o <= 16'h0000;
        10'h2b5: pm_insn_o <= 16'h0000;
        10'h2b6: pm_insn_o <= 16'h0000;
        10'h2b7: pm_insn_o <= 16'h0000;
        10'h2b8: pm_insn_o <= 16'h0000;
        10'h2b9: pm_insn_o <= 16'h0000;
        10'h2ba: pm_insn_o <= 16'h0000;
        10'h2bb: pm_insn_o <= 16'h0000;
        10'h2bc: pm_insn_o <= 16'h0000;
        10'h2bd: pm_insn_o <= 16'h0000;
        10'h2be: pm_insn_o <= 16'h0000;
        10'h2bf: pm_insn_o <= 16'h0000;
        10'h2c0: pm_insn_o <= 16'h0000;
        10'h2c1: pm_insn_o <= 16'h0000;
        10'h2c2: pm_insn_o <= 16'h0000;
        10'h2c3: pm_insn_o <= 16'h0000;
        10'h2c4: pm_insn_o <= 16'h0000;
        10'h2c5: pm_insn_o <= 16'h0000;
        10'h2c6: pm_insn_o <= 16'h0000;
        10'h2c7: pm_insn_o <= 16'h0000;
        10'h2c8: pm_insn_o <= 16'h0000;
        10'h2c9: pm_insn_o <= 16'h0000;
        10'h2ca: pm_insn_o <= 16'h0000;
        10'h2cb: pm_insn_o <= 16'h0000;
        10'h2cc: pm_insn_o <= 16'h0000;
        10'h2cd: pm_insn_o <= 16'h0000;
        10'h2ce: pm_insn_o <= 16'h0000;
        10'h2cf: pm_insn_o <= 16'h0000;
        10'h2d0: pm_insn_o <= 16'h0000;
        10'h2d1: pm_insn_o <= 16'h0000;
        10'h2d2: pm_insn_o <= 16'h0000;
        10'h2d3: pm_insn_o <= 16'h0000;
        10'h2d4: pm_insn_o <= 16'h0000;
        10'h2d5: pm_insn_o <= 16'h0000;
        10'h2d6: pm_insn_o <= 16'h0000;
        10'h2d7: pm_insn_o <= 16'h0000;
        10'h2d8: pm_insn_o <= 16'h0000;
        10'h2d9: pm_insn_o <= 16'h0000;
        10'h2da: pm_insn_o <= 16'h0000;
        10'h2db: pm_insn_o <= 16'h0000;
        10'h2dc: pm_insn_o <= 16'h0000;
        10'h2dd: pm_insn_o <= 16'h0000;
        10'h2de: pm_insn_o <= 16'h0000;
        10'h2df: pm_insn_o <= 16'h0000;
        10'h2e0: pm_insn_o <= 16'h0000;
        10'h2e1: pm_insn_o <= 16'h0000;
        10'h2e2: pm_insn_o <= 16'h0000;
        10'h2e3: pm_insn_o <= 16'h0000;
        10'h2e4: pm_insn_o <= 16'h0000;
        10'h2e5: pm_insn_o <= 16'h0000;
        10'h2e6: pm_insn_o <= 16'h0000;
        10'h2e7: pm_insn_o <= 16'h0000;
        10'h2e8: pm_insn_o <= 16'h0000;
        10'h2e9: pm_insn_o <= 16'h0000;
        10'h2ea: pm_insn_o <= 16'h0000;
        10'h2eb: pm_insn_o <= 16'h0000;
        10'h2ec: pm_insn_o <= 16'h0000;
        10'h2ed: pm_insn_o <= 16'h0000;
        10'h2ee: pm_insn_o <= 16'h0000;
        10'h2ef: pm_insn_o <= 16'h0000;
        10'h2f0: pm_insn_o <= 16'h0000;
        10'h2f1: pm_insn_o <= 16'h0000;
        10'h2f2: pm_insn_o <= 16'h0000;
        10'h2f3: pm_insn_o <= 16'h0000;
        10'h2f4: pm_insn_o <= 16'h0000;
        10'h2f5: pm_insn_o <= 16'h0000;
        10'h2f6: pm_insn_o <= 16'h0000;
        10'h2f7: pm_insn_o <= 16'h0000;
        10'h2f8: pm_insn_o <= 16'h0000;
        10'h2f9: pm_insn_o <= 16'h0000;
        10'h2fa: pm_insn_o <= 16'h0000;
        10'h2fb: pm_insn_o <= 16'h0000;
        10'h2fc: pm_insn_o <= 16'h0000;
        10'h2fd: pm_insn_o <= 16'h0000;
        10'h2fe: pm_insn_o <= 16'h0000;
        10'h2ff: pm_insn_o <= 16'h0000;
        10'h300: pm_insn_o <= 16'h0d0a; // 	dw	0x0d0a
        10'h301: pm_insn_o <= 16'h4145; // 	dw	0x4145
        10'h302: pm_insn_o <= 16'h0000; // 	dw	0x0000
        10'h303: pm_insn_o <= 16'h0000;
        10'h304: pm_insn_o <= 16'h0000;
        10'h305: pm_insn_o <= 16'h0000;
        10'h306: pm_insn_o <= 16'h0000;
        10'h307: pm_insn_o <= 16'h0000;
        10'h308: pm_insn_o <= 16'h0000;
        10'h309: pm_insn_o <= 16'h0000;
        10'h30a: pm_insn_o <= 16'h0000;
        10'h30b: pm_insn_o <= 16'h0000;
        10'h30c: pm_insn_o <= 16'h0000;
        10'h30d: pm_insn_o <= 16'h0000;
        10'h30e: pm_insn_o <= 16'h0000;
        10'h30f: pm_insn_o <= 16'h0000;
        10'h310: pm_insn_o <= 16'h0000;
        10'h311: pm_insn_o <= 16'h0000;
        10'h312: pm_insn_o <= 16'h0000;
        10'h313: pm_insn_o <= 16'h0000;
        10'h314: pm_insn_o <= 16'h0000;
        10'h315: pm_insn_o <= 16'h0000;
        10'h316: pm_insn_o <= 16'h0000;
        10'h317: pm_insn_o <= 16'h0000;
        10'h318: pm_insn_o <= 16'h0000;
        10'h319: pm_insn_o <= 16'h0000;
        10'h31a: pm_insn_o <= 16'h0000;
        10'h31b: pm_insn_o <= 16'h0000;
        10'h31c: pm_insn_o <= 16'h0000;
        10'h31d: pm_insn_o <= 16'h0000;
        10'h31e: pm_insn_o <= 16'h0000;
        10'h31f: pm_insn_o <= 16'h0000;
        10'h320: pm_insn_o <= 16'h0000;
        10'h321: pm_insn_o <= 16'h0000;
        10'h322: pm_insn_o <= 16'h0000;
        10'h323: pm_insn_o <= 16'h0000;
        10'h324: pm_insn_o <= 16'h0000;
        10'h325: pm_insn_o <= 16'h0000;
        10'h326: pm_insn_o <= 16'h0000;
        10'h327: pm_insn_o <= 16'h0000;
        10'h328: pm_insn_o <= 16'h0000;
        10'h329: pm_insn_o <= 16'h0000;
        10'h32a: pm_insn_o <= 16'h0000;
        10'h32b: pm_insn_o <= 16'h0000;
        10'h32c: pm_insn_o <= 16'h0000;
        10'h32d: pm_insn_o <= 16'h0000;
        10'h32e: pm_insn_o <= 16'h0000;
        10'h32f: pm_insn_o <= 16'h0000;
        10'h330: pm_insn_o <= 16'h0000;
        10'h331: pm_insn_o <= 16'h0000;
        10'h332: pm_insn_o <= 16'h0000;
        10'h333: pm_insn_o <= 16'h0000;
        10'h334: pm_insn_o <= 16'h0000;
        10'h335: pm_insn_o <= 16'h0000;
        10'h336: pm_insn_o <= 16'h0000;
        10'h337: pm_insn_o <= 16'h0000;
        10'h338: pm_insn_o <= 16'h0000;
        10'h339: pm_insn_o <= 16'h0000;
        10'h33a: pm_insn_o <= 16'h0000;
        10'h33b: pm_insn_o <= 16'h0000;
        10'h33c: pm_insn_o <= 16'h0000;
        10'h33d: pm_insn_o <= 16'h0000;
        10'h33e: pm_insn_o <= 16'h0000;
        10'h33f: pm_insn_o <= 16'h0000;
        10'h340: pm_insn_o <= 16'h0000;
        10'h341: pm_insn_o <= 16'h0000;
        10'h342: pm_insn_o <= 16'h0000;
        10'h343: pm_insn_o <= 16'h0000;
        10'h344: pm_insn_o <= 16'h0000;
        10'h345: pm_insn_o <= 16'h0000;
        10'h346: pm_insn_o <= 16'h0000;
        10'h347: pm_insn_o <= 16'h0000;
        10'h348: pm_insn_o <= 16'h0000;
        10'h349: pm_insn_o <= 16'h0000;
        10'h34a: pm_insn_o <= 16'h0000;
        10'h34b: pm_insn_o <= 16'h0000;
        10'h34c: pm_insn_o <= 16'h0000;
        10'h34d: pm_insn_o <= 16'h0000;
        10'h34e: pm_insn_o <= 16'h0000;
        10'h34f: pm_insn_o <= 16'h0000;
        10'h350: pm_insn_o <= 16'h0000;
        10'h351: pm_insn_o <= 16'h0000;
        10'h352: pm_insn_o <= 16'h0000;
        10'h353: pm_insn_o <= 16'h0000;
        10'h354: pm_insn_o <= 16'h0000;
        10'h355: pm_insn_o <= 16'h0000;
        10'h356: pm_insn_o <= 16'h0000;
        10'h357: pm_insn_o <= 16'h0000;
        10'h358: pm_insn_o <= 16'h0000;
        10'h359: pm_insn_o <= 16'h0000;
        10'h35a: pm_insn_o <= 16'h0000;
        10'h35b: pm_insn_o <= 16'h0000;
        10'h35c: pm_insn_o <= 16'h0000;
        10'h35d: pm_insn_o <= 16'h0000;
        10'h35e: pm_insn_o <= 16'h0000;
        10'h35f: pm_insn_o <= 16'h0000;
        10'h360: pm_insn_o <= 16'h0000;
        10'h361: pm_insn_o <= 16'h0000;
        10'h362: pm_insn_o <= 16'h0000;
        10'h363: pm_insn_o <= 16'h0000;
        10'h364: pm_insn_o <= 16'h0000;
        10'h365: pm_insn_o <= 16'h0000;
        10'h366: pm_insn_o <= 16'h0000;
        10'h367: pm_insn_o <= 16'h0000;
        10'h368: pm_insn_o <= 16'h0000;
        10'h369: pm_insn_o <= 16'h0000;
        10'h36a: pm_insn_o <= 16'h0000;
        10'h36b: pm_insn_o <= 16'h0000;
        10'h36c: pm_insn_o <= 16'h0000;
        10'h36d: pm_insn_o <= 16'h0000;
        10'h36e: pm_insn_o <= 16'h0000;
        10'h36f: pm_insn_o <= 16'h0000;
        10'h370: pm_insn_o <= 16'h0000;
        10'h371: pm_insn_o <= 16'h0000;
        10'h372: pm_insn_o <= 16'h0000;
        10'h373: pm_insn_o <= 16'h0000;
        10'h374: pm_insn_o <= 16'h0000;
        10'h375: pm_insn_o <= 16'h0000;
        10'h376: pm_insn_o <= 16'h0000;
        10'h377: pm_insn_o <= 16'h0000;
        10'h378: pm_insn_o <= 16'h0000;
        10'h379: pm_insn_o <= 16'h0000;
        10'h37a: pm_insn_o <= 16'h0000;
        10'h37b: pm_insn_o <= 16'h0000;
        10'h37c: pm_insn_o <= 16'h0000;
        10'h37d: pm_insn_o <= 16'h0000;
        10'h37e: pm_insn_o <= 16'h0000;
        10'h37f: pm_insn_o <= 16'h0000;
        10'h380: pm_insn_o <= 16'h0000;
        10'h381: pm_insn_o <= 16'h0000;
        10'h382: pm_insn_o <= 16'h0000;
        10'h383: pm_insn_o <= 16'h0000;
        10'h384: pm_insn_o <= 16'h0000;
        10'h385: pm_insn_o <= 16'h0000;
        10'h386: pm_insn_o <= 16'h0000;
        10'h387: pm_insn_o <= 16'h0000;
        10'h388: pm_insn_o <= 16'h0000;
        10'h389: pm_insn_o <= 16'h0000;
        10'h38a: pm_insn_o <= 16'h0000;
        10'h38b: pm_insn_o <= 16'h0000;
        10'h38c: pm_insn_o <= 16'h0000;
        10'h38d: pm_insn_o <= 16'h0000;
        10'h38e: pm_insn_o <= 16'h0000;
        10'h38f: pm_insn_o <= 16'h0000;
        10'h390: pm_insn_o <= 16'h0000;
        10'h391: pm_insn_o <= 16'h0000;
        10'h392: pm_insn_o <= 16'h0000;
        10'h393: pm_insn_o <= 16'h0000;
        10'h394: pm_insn_o <= 16'h0000;
        10'h395: pm_insn_o <= 16'h0000;
        10'h396: pm_insn_o <= 16'h0000;
        10'h397: pm_insn_o <= 16'h0000;
        10'h398: pm_insn_o <= 16'h0000;
        10'h399: pm_insn_o <= 16'h0000;
        10'h39a: pm_insn_o <= 16'h0000;
        10'h39b: pm_insn_o <= 16'h0000;
        10'h39c: pm_insn_o <= 16'h0000;
        10'h39d: pm_insn_o <= 16'h0000;
        10'h39e: pm_insn_o <= 16'h0000;
        10'h39f: pm_insn_o <= 16'h0000;
        10'h3a0: pm_insn_o <= 16'h0000;
        10'h3a1: pm_insn_o <= 16'h0000;
        10'h3a2: pm_insn_o <= 16'h0000;
        10'h3a3: pm_insn_o <= 16'h0000;
        10'h3a4: pm_insn_o <= 16'h0000;
        10'h3a5: pm_insn_o <= 16'h0000;
        10'h3a6: pm_insn_o <= 16'h0000;
        10'h3a7: pm_insn_o <= 16'h0000;
        10'h3a8: pm_insn_o <= 16'h0000;
        10'h3a9: pm_insn_o <= 16'h0000;
        10'h3aa: pm_insn_o <= 16'h0000;
        10'h3ab: pm_insn_o <= 16'h0000;
        10'h3ac: pm_insn_o <= 16'h0000;
        10'h3ad: pm_insn_o <= 16'h0000;
        10'h3ae: pm_insn_o <= 16'h0000;
        10'h3af: pm_insn_o <= 16'h0000;
        10'h3b0: pm_insn_o <= 16'h0000;
        10'h3b1: pm_insn_o <= 16'h0000;
        10'h3b2: pm_insn_o <= 16'h0000;
        10'h3b3: pm_insn_o <= 16'h0000;
        10'h3b4: pm_insn_o <= 16'h0000;
        10'h3b5: pm_insn_o <= 16'h0000;
        10'h3b6: pm_insn_o <= 16'h0000;
        10'h3b7: pm_insn_o <= 16'h0000;
        10'h3b8: pm_insn_o <= 16'h0000;
        10'h3b9: pm_insn_o <= 16'h0000;
        10'h3ba: pm_insn_o <= 16'h0000;
        10'h3bb: pm_insn_o <= 16'h0000;
        10'h3bc: pm_insn_o <= 16'h0000;
        10'h3bd: pm_insn_o <= 16'h0000;
        10'h3be: pm_insn_o <= 16'h0000;
        10'h3bf: pm_insn_o <= 16'h0000;
        10'h3c0: pm_insn_o <= 16'h0000;
        10'h3c1: pm_insn_o <= 16'h0000;
        10'h3c2: pm_insn_o <= 16'h0000;
        10'h3c3: pm_insn_o <= 16'h0000;
        10'h3c4: pm_insn_o <= 16'h0000;
        10'h3c5: pm_insn_o <= 16'h0000;
        10'h3c6: pm_insn_o <= 16'h0000;
        10'h3c7: pm_insn_o <= 16'h0000;
        10'h3c8: pm_insn_o <= 16'h0000;
        10'h3c9: pm_insn_o <= 16'h0000;
        10'h3ca: pm_insn_o <= 16'h0000;
        10'h3cb: pm_insn_o <= 16'h0000;
        10'h3cc: pm_insn_o <= 16'h0000;
        10'h3cd: pm_insn_o <= 16'h0000;
        10'h3ce: pm_insn_o <= 16'h0000;
        10'h3cf: pm_insn_o <= 16'h0000;
        10'h3d0: pm_insn_o <= 16'h0000;
        10'h3d1: pm_insn_o <= 16'h0000;
        10'h3d2: pm_insn_o <= 16'h0000;
        10'h3d3: pm_insn_o <= 16'h0000;
        10'h3d4: pm_insn_o <= 16'h0000;
        10'h3d5: pm_insn_o <= 16'h0000;
        10'h3d6: pm_insn_o <= 16'h0000;
        10'h3d7: pm_insn_o <= 16'h0000;
        10'h3d8: pm_insn_o <= 16'h0000;
        10'h3d9: pm_insn_o <= 16'h0000;
        10'h3da: pm_insn_o <= 16'h0000;
        10'h3db: pm_insn_o <= 16'h0000;
        10'h3dc: pm_insn_o <= 16'h0000;
        10'h3dd: pm_insn_o <= 16'h0000;
        10'h3de: pm_insn_o <= 16'h0000;
        10'h3df: pm_insn_o <= 16'h0000;
        10'h3e0: pm_insn_o <= 16'h0000;
        10'h3e1: pm_insn_o <= 16'h0000;
        10'h3e2: pm_insn_o <= 16'h0000;
        10'h3e3: pm_insn_o <= 16'h0000;
        10'h3e4: pm_insn_o <= 16'h0000;
        10'h3e5: pm_insn_o <= 16'h0000;
        10'h3e6: pm_insn_o <= 16'h0000;
        10'h3e7: pm_insn_o <= 16'h0000;
        10'h3e8: pm_insn_o <= 16'h0000;
        10'h3e9: pm_insn_o <= 16'h0000;
        10'h3ea: pm_insn_o <= 16'h0000;
        10'h3eb: pm_insn_o <= 16'h0000;
        10'h3ec: pm_insn_o <= 16'h0000;
        10'h3ed: pm_insn_o <= 16'h0000;
        10'h3ee: pm_insn_o <= 16'h0000;
        10'h3ef: pm_insn_o <= 16'h0000;
        10'h3f0: pm_insn_o <= 16'h0000;
        10'h3f1: pm_insn_o <= 16'h0000;
        10'h3f2: pm_insn_o <= 16'h0000;
        10'h3f3: pm_insn_o <= 16'h0000;
        10'h3f4: pm_insn_o <= 16'h0000;
        10'h3f5: pm_insn_o <= 16'h0000;
        10'h3f6: pm_insn_o <= 16'h0000;
        10'h3f7: pm_insn_o <= 16'h0000;
        10'h3f8: pm_insn_o <= 16'h0000;
        10'h3f9: pm_insn_o <= 16'h0000;
        10'h3fa: pm_insn_o <= 16'h0000;
        10'h3fb: pm_insn_o <= 16'h0000;
        10'h3fc: pm_insn_o <= 16'h0000;
        10'h3fd: pm_insn_o <= 16'h0000;
        10'h3fe: pm_insn_o <= 16'h0000;
        10'h3ff: pm_insn_o <= 16'hab54; // 	dw	0xab54		; Just a check intended for tools that automatically poke around inside this memory
        default: pm_insn_o <= 16'h0000;
      endcase // case(pm_addr_i)

endmodule // serial_wb_program
